module turbo_test();

reg[6143:0] in;
reg[6143:0] out;
reg[6143:0] expected_out;

integer counter, counter_rev;
reg start_rec;
reg start_send;

//inputs
reg clk, reset, vld_crc, rdy_out, cbs;
reg [7:0] data_in_rev;
reg [7:0] data_in;

//outputs
wire rdy_crc, vld_out, last_byte;
wire [7:0] data_out;

string correct;

initial 
begin

$display("starting simulation");
$display("counter | reset | vld_crc | where_in_block | data_in");

in <= 6144'b010101001101000101111110101101110000010010011011101111110010100110111011001011100110101000111010001100000011100100110110010100001010010011011111111111111110110111001001100101001111111111100100010101110101110101101101000101101000101110010011111000011000111111111111111110010000101011010011101101010100011001111010001001011001111110101001110101100100101011011011011111001010000010000100011000101010111000010101100011110000101101111110000100000110001111111101110101101111101011010100000000100010001111100101101011110010001101010100011100100110000000000001011101100001010111110101010011101000010001001101111000010011001100111101111010011000000100100110101111101110111100111000110111010000100110000110000110010001000110110100101111000110110111000001110110101101101001010111111100000101100011010110010001000001111101111101100010011000110110101110110111100100011000111001011101000110100000001010100101011010001011010011000011100101011101010101010100001011000110111100111001111011101101111010001110100110001010010000111010011010111110001001000010100111001100000001111111101110110111000011001100110111001101111010010101011000001110000101011100000011101000001000000000110000011000011100000010111101100010000011001000010100000010100010100101111011000000110111110001100010011100101101110001100110100111011110100001000000110100110110000001001000101000011011110111111110001110100111000011101100001001001010000010100000011000100000010010011110010011111100101100111101010101110000110010011000111110010111010011011010100100010101010110010010010111000101011100100101000101101010111011011000011111101001100111010110000011111011100010001011111100000000101100101001111111001001100010001011001111010101001100100110110010011010111110110100101010111110001011101001110101001100011100010111001110000111110000101111001100001011111010110001000110111101010010001111000010101110110111000101101100000000100011111010110010100101101000111010001001011100010110011101000110100101110011101100011000111001110000110110111100110100000110000101011000000000011110111101000110110111010111000111101001010001101111001010100001100001011101000011001101001111101101101000110101101110100111011101110001110010000110011011111101001100010111100010100000001000110011100100011001101111100000100000110100101010100000010010100110110000000011011010010000001010110010000110000010110000101100110001110000011001001100010001011100011100100010001100100011011010011111101110011010111110111100000111010111100001010100100100111011000011011000100111101001110011110100000010100101011000010101110010111010100011110111101001011111011111100011001100101000100110110110100100011101101100011010100100000001000101000111110111000000100001011110100100010011111001100010110001001110011100110000110101101110011110110110011111110001011100100010001011011110101101011111000001001110011101111000001011010010010011101011110000101100111011100010110111011010111101101111111101100001000110100111000100001011010011010110100101111000011000000000001000110000101010111110000001110010100100010111101100111101010010101001001110101111011111011000011011100001011111010001000110000001101101111110010000100111100100001000110101111100101101101100111001101011110001100100101010001111110101001110101110100010101111111100010100011011011101101100100011001111110000010111001101111010101011110010010001010100001011110011100110101110110011011001000011110010010111111011111000000010001001000000001110000111001111100101111110011110010011010001110100111111011100111110101101011000101101101000011010100000011100100110100101111011111010011010000101001100110110000111000010010000100011100010011100000100010010010111000100010111111011111000110101100101000110111011100110111100010101111001111110111100110101010101101000011001101100111001110010010110000011011100010111110010010110000101100000011110100100011011100010000101100001010011100101011011010011101111001011001000101010010110000010100100110000011111111000001010000001110001110001110011010001101111010100001001100000000000100001010010100010100101000100010000110100101011110111101001110101110111100111101001100111010000101001011001000001000101011101010111000011011010110100111110001100011000101010000010101010000011011001001000100000010100100100111000000010011001111110001000010010110110110100100100011001001100100010100100000001111011101110010111000001100110111010010011001000111001111001110111000110110110001011111000100111100111100111111010000100101110000011111001011001010001101101110011100111110101001010111110101010111011111001010000011010011011010011111010000001000011001001111101010100100111010111100000001010110001011011010000010011000011101100111000110100010100001100100110110010100100110001100011110010101111001110101101001100011000100101100001011101110000101010100111001100100011001000100110001001111011010100010111111111101011010111100000001100010010010001101001111011001011110111010000000001010111010001001010001101001010101100110110001101010001111111110000110110100101010110100000010010011101000111011111010100000111101100101101101001101110100100001101010100110000011001100100101001100110010010001010111110101111100100101111110000001101100001011010100011111100001110011001100000111111111111010010111010001111001111100010010011100110011001101101111110011001001110100110000001011100110101000110001011101110011111000011001001010100000111001000101100000010001010000011111011100001000001011001100111110010110011001101100010001011111110011001110010100011011100101001011010000101010010100111100110000000011000111010110100100110000011011101000000011110100110110011111001110011010011001000110011100010110101100101101010010010011101001110011000111100001100011001000010010010010000000100001010110101101101000000111101010110111101001011001000001010001101111001010110000001100110010111101111010100100110000010000001111110101010011001101111111011101111010001110010100111000001011011000000010111101111011000000000010101111111110100011101101101001011001001110111111000000100010111100001100000001011110101000110000001111001000011010000000101111100110011001101111111101010001001101101011111111001000000000101111111001001100000101010100001111101011010101010111110011111101000110000010110001101100111011001;
expected_out <= 6144'b010000110010100111101101110011011100010001001011100100001101111100101000110011110010111011010010100101111001011110100001110000010110010001101010110100101011101011001101000000011100110110011001110001011100000001001101001001011000111000101100000100001011111110110101101001110111101011010000001001101100000001111110001011001100101111111011000101101111000001111100000001101010101010000000110010100111000111110101111101101011001100011000100101010110001000010100001110010000111100001110111000101000001011001001001101000101100000110011010110000101110100111101010111111100010110001000110101111101111100000100011101101010110001111011110111011011010100100101100011101011000001101110100110110000000010001110010000101111011000011111101100111100001100111011011110000100111010110011000111110101101001001000111100000110000000001110010001001011101100100011101000011000111101110001100101100110111000110101000101110000000011101111110000110110111111110111110000010110010010001001001001001110010100110111101101010110100101101001001011010001001011011101010000001000010001011001100101001110100111010110011101101100110001101110100000010001001010010110010000000100011010011000011001000101100110001100000110010010000110111010100000100000110110011101111100110000111000100101110001000111101111000010111000111011111111100010011110000110110100101101101111100000110100100110001100110100010111110110010011000001100110010011010010100010111010100011010010010110011110000000101101110111101100011111010101111100011110101001110000001101011000010000110011000011110001110110011000111110110000001011101000101111110000100001001110101111101111000101111010001110111110111111010010000010000001110001001101000010011000101010010100001000000010010011101110100111111111000010011110010001110000010000010110100010101101001011101111100111011010110011000001111011000011100000001011000010110101110111111011100010001100110001100011111101100110011100001001000011010010000000011100101000011000011011001101111000001100100010000001010101001111011001110011111001100010111011010111111100001010100111011001011010000101001000000011110001011111110011101100011101100110011111111001000100000000100111001011111001010100001001110111100000011010010100010110001110011011011100111100011000100011111000010001001001111101010000101011000010110110101100101001010100001010000111111100000000110010011111110011110110001110111100000010101100100100101110100101000101111010111010010111001000100111001100001000100000011111110010000011010111001100111111100001000011000101101000111001010110000000001011100010010000010010011111110010011111010011110110011110001001101100100100011010011101111101111000011101000100001010100011101000000100110000101110011110111101101011110001011010100110100011001101011011100111001101110010100111001100101101111000111011011100011001100001110100001111001110001111100101001011011101001111001000100111010011111011110010110011110110101111010111111001100110101101100010100111010110001111110001110010001110000010111010101000100100011011010111011100010110000001110111100010010010010111111110110011111000100000110001110000001110101111010110001101101100000110110001010011001101001101110110001100001110100110100011001011111110011110001101110101001001111001101010100100100100100100000001001000010011111101001101100001000001100000000010011010111001011101000010110100101001110000100101011010011110001111110001100010000000001000001101100110101111000101101010111011000100100100011100000011000011000001100000000100011101010110110110001010001001011011100011111001001100100000101100010101110111100101001111110010111110110010111011111110111001000101100110101111000010110111111010001111001001010111010111000110001001100010101001010000000111011010010011111010001101100100111001101110110100111001111001000011000110010111100100001001101010011000100001101001100111110110110110010011001000111100110111010001101101101101110111010010001110010001011011000000100000000100000100011010101101111011100000010001010100011100101111001010001001010101110110101000100001111101100100000101111110110110111010101101011000110001101110011010110101001101000010011111010011101111111110001010110000000010011011010011001001001100100000001100000111111110011000101000101011001111100010100000110100001110001011011011000010001011111010011011011110110011010111001100010000111001100000011110111110100001000001100010111000100000010010110010001100100100011101100000110111010000111100010011110111011111101010110100100101011000010110110011111100011110000010111001000011001101001101100011100110111111001011001001010011111100011010010101110101111011010111000110011000000001001100000100011010111100000001000001100111011101001111100111101101001111111000110001110100010100100011011101110111000010000001111111011101001101101111001111101001101101110100010101001101110111110000111011000001011100110110100010010000111111111100000111000111001101001110011001000010100001100001011101010001101010010100010010000110011110010011110100000111110000110010001100111110101100000010011110011011011101001101100010001010000001100110111011011111011001101111011111100000011001110101100101111001110010111010101010110100001011001010110111101011001001111000101110010001010000000101101001000100100010111011011000001110101001010101011111110100101101001010111101010101110101110010110101101100001111101111011001110010101000001110000011100111011001101111000110000011001101010001111110010001010110110001011000000001100100111100011001100011111100011111111111010110011000001101011011010010010101101011111110001100011110100100010010111010100101111101110101101000000000101001000011101010010111101000100011010111011100111010110001100110111011010110101001100100111111000011110000011100001100010011101010001101101101000100101100100000010101000100111010111111111001001000101011000011110001100110100000010010011101101101100001000000111000110110111100110000101101001000000001101000100100001000100111110011110101011101000111010000101111100100011010100101100100101001010001110100110101110000100010011001000111011100000101101100010001001100100100101110111110110010100010100111101110000111100111011110000010111111101010101001101001110000101011100111001110111011111110101100010000011111101011110100110000;
reset <= 1'b1;
vld_crc <= 1'b0;
rdy_out <= 1'b0;
clk <= 1'b0;
start_rec <= 1'b0;
start_send <= 1'b0;
cbs <= 1'b1;

counter <= 0;

data_in <= 8'd0;
data_in_rev <= 8'd0;


end

always
begin
#10 clk <= ~clk;
end

//inital reset and setup
always
begin
//reset
@(posedge clk)
@(posedge clk)
@(posedge clk)
//end reset and assert vld_crc
@(negedge clk) begin
 reset <= 1'b0;
 vld_crc <= 1'b1;
end
@(posedge rdy_crc) begin
 rdy_out <= 1'b1;
 counter <= 0;
end

//wait until we get vld_out
@(posedge vld_out) begin
 vld_crc <= 1'b0;
end

@(posedge clk) begin
	counter <= 0;
end

#3000
$stop;
end

always @(negedge clk)
begin
	if(rdy_crc) begin
		counter_rev = (6144 - counter) - 8;
		counter = counter + 8;	
	end
	if(vld_out) begin
		counter_rev = (6144 - counter) - 8;
		counter = counter + 8;
	end
	// if recieving
	if(rdy_crc) begin
		data_in = in[counter_rev +: 8];
//		data_in[0] <= data_in_rev[7];
//		data_in[1] <= data_in_rev[6];
//		data_in[2] <= data_in_rev[5];
//		data_in[3] <= data_in_rev[4];
//		data_in[4] <= data_in_rev[3];
//		data_in[5] <= data_in_rev[2];
//		data_in[6] <= data_in_rev[1];
//		data_in[7] <= data_in_rev[0];
	end
	//if sending
	if(vld_out) begin
		out[counter_rev +: 8] = data_out;
		if(data_out == expected_out[counter_rev +: 8])
		begin
			correct = "TRUE";
		end
		else 
		begin
			correct = "FALSE";
		end
	end
	
	
end

always @(posedge clk) begin
	$display("count: %0d | vld_crc: %b | rdy_crc: %b | vld_out: %b | last_byte: %b | data_in: %b | data_out: %b | expected: %b | correct: %s", counter_rev, vld_crc, rdy_crc, vld_out, last_byte, data_in, data_out, expected_out[counter_rev +: 8], correct);
end

interleaver dut(clk, reset, vld_crc, rdy_out, cbs, data_in, rdy_crc, vld_out, last_byte, data_out);


endmodule
