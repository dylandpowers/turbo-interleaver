module turbo_test();

reg[1055:0] in;
reg[1055:0] out;
reg[1055:0] expected_out;

integer counter, counter_rev;
reg start_rec;
reg start_send;

//inputs
reg clk, reset, vld_crc, rdy_out, cbs;
reg [7:0] data_in_rev;
reg [7:0] data_in;

//outputs
wire rdy_crc, vld_out, last_byte;
wire [7:0] data_out;

string correct;

initial 
begin

$display("starting simulation");
$display("counter | reset | vld_crc | where_in_block | data_in");

in <= 1056'b010011010101110101100111100000011111001001010101100011011101011000101001111001010110010001001000011100100001010001110000010110100011101011100110001001001110011000000000100110000100110111101000001101001011100101011011100100111100011111001001000100010000011111011110001001011011001001010000101010101110011000110110000100110111010100000011101010010111000111111101111100000010110101101101010110101101001011000101011001011101111111000010000100001011011010100100000111101010101000010101001111110100100100011000100011100011111011100010110011001101000011000010111011011011001111000110100010010111111011101010010111010101010001101001010111100101011001111010101100100111111010110001001110001111000000110010110111011011100001100000001010010110111010110110001100011100111011110100000100001011000101010001111011010000100111100011011101111110001010001110001111011000110011111001101010110011111110101110001111000100111110110110101001111110011011011010110111100011010100100001111101001000010101110100000000010101101011011010101001000011110010101110001010110000001100111110;
expected_out <= 1056'b001010011100110111011110001101011110001111110010000110110010101111000010101011010101100110101001111010110011011111000010010111110010101011010111110100010001001101111101000000011100000101010000000100111101001100110111110000100001101111101001111000110011010101000100011100101100110110001010000100111100100100110111111011110100001110110110011111011111001111000100001000000000000010111010010111010001001010111010010001011111110100111101110000110101000011101111111001010011000100001111000110001010001100011000010111101011000011101110111010011111101000001100110011000101000010110010101010101011110111111110110001001011101011011011111001011010011000111000010101111111110000101110110111001001111000100010101000011110100100011000011001011100010001110000011000000111110100010000001101011111101001101000111111111001100100100000001011100101011011111001110110100100101011111010101011010110000101010001010011001010111101100100001101001111010000001011101001010001001100100001011000000110010010100111001100011011001100001110010101010111001000101011101001000001110011010010;
reset <= 1'b1;
vld_crc <= 1'b0;
rdy_out <= 1'b0;
clk <= 1'b0;
start_rec <= 1'b0;
start_send <= 1'b0;
cbs <= 1'b0;

counter <= 0;

data_in <= 8'd0;
data_in_rev <= 8'd0;


end

always
begin
#10 clk <= ~clk;
end

//inital reset and setup
always
begin
//reset
@(posedge clk)
@(posedge clk)
@(posedge clk)
//end reset and assert vld_crc
@(negedge clk) begin
 reset <= 1'b0;
 vld_crc <= 1'b1;
end
@(posedge rdy_crc) begin
 rdy_out <= 1'b1;
 counter <= 0;
end

//wait until we get vld_out
@(posedge vld_out) begin
 vld_crc <= 1'b0;
end

@(posedge clk) begin
	counter <= 0;
end

#3000
$stop;
end

always @(negedge clk)
begin
	if(rdy_crc) begin
		counter_rev = (1056 - counter) - 8;
		counter = counter + 8;	
	end
	if(vld_out) begin
		counter_rev = (1056 - counter) - 8;
		counter = counter + 8;
	end
	// if recieving
	if(rdy_crc) begin
		data_in = in[counter_rev +: 8];
//		data_in[0] <= data_in_rev[7];
//		data_in[1] <= data_in_rev[6];
//		data_in[2] <= data_in_rev[5];
//		data_in[3] <= data_in_rev[4];
//		data_in[4] <= data_in_rev[3];
//		data_in[5] <= data_in_rev[2];
//		data_in[6] <= data_in_rev[1];
//		data_in[7] <= data_in_rev[0];
	end
	//if sending
	if(vld_out) begin
		out[counter_rev +: 8] = data_out;
		if(data_out == expected_out[counter_rev +: 8])
		begin
			correct = "TRUE";
		end
		else 
		begin
			correct = "FALSE";
		end
	end
	
	
end

always @(posedge clk) begin
	$display("count: %0d | vld_crc: %b | rdy_crc: %b | vld_out: %b | last_byte: %b | data_in: %b | data_out: %b | expected: %b | correct: %s", counter_rev, vld_crc, rdy_crc, vld_out, last_byte, data_in, data_out, expected_out[counter_rev +: 8], correct);
end

interleaver dut(clk, reset, vld_crc, rdy_out, cbs, data_in, rdy_crc, vld_out, last_byte, data_out);


endmodule
