module turbo_test();

reg[1055:0] in;
reg[1055:0] out;
reg[1055:0] expected_out;

integer counter;
reg[31:0] where_in_block;
reg[31:0] where_in_block7;
reg start_rec;
reg start_send;

//inputs
reg clk, reset, vld_crc, rdy_out, cbs;
reg[7:0] data_in;

//outputs
wire rdy_crc, vld_out;
wire[7:0] data_out;

string correct;

initial 
begin

	$display("starting simulation");
	$display("counter | reset | vld_crc | where_in_block | data_in");
	
	in <= 1056'b111011000111110000011110000110000101111100001010110100011111000111100010001011010010000100100100100001000111100100001000110110100101001110111100100100100111101001101111111101111011100100011111010001111100100111110001101101010011110101010110101110001011000111100111101110000001100110101100011001011000011111010111111111110011110011101111110110010000111010110100110001100011100001111011001110110011011010000101001101010010010111011101110101010110001110101010111110000110100011100100000010101000110110110010010000110010000110100010110001111010011010110000000011010110100000000011100001101111011010011010110000110111110011011110111111110000011011100110101110011100101100100110010001111000000101001101011100010000111111000111101111101001111001111000001011010000100111110100001111011111000011011000010111100101000101111011101010100111001110001010010110011111001110110100010000111110101010100010001111111101010110000110011101010011010110000111001011111010101101110011100011011111110101100111001000011100111000110110110110111001000010000011100010111011101011101011;
	expected_out <= 1056'b100101101100111001011111000000001100111011101111111101100001011000110110111001101100111000100101101101111101011110110010011011001101000010101000100101001010001100010101011110001000101110101000111011000100001000100010010100111111111111011000001001001011000001010101101111101010100111000000001111100101110110011000011101110110101011010110100101110100011001111000011100100010100111101000010001011111000001100110100101010001001011001101111011100111101001100110100111101000100000010110011111011001100110110111101110111101111100001000111010110000101100000100011001010010011101110101011101011011100100101100010101001111000010111000110110010100000000011001100001111010111111011011001000110111101100110110101111101111011010011111101010011111011010101100110111010010100010111101000010001010001011101101000001011110101100001101111000111001111101011101001111010110111100111111110000000100110010101111111011101011001010111110110111001000001011011011011111011000101001100011001000001110001100101000010101101111101101010001111001110100010101110111111100101000010101100001;
	cbs <= 1'b0;
	reset <= 1'b1;
	vld_crc <= 1'b0;
	rdy_out <= 1'b0;
	clk <= 1'b0;
	
	counter <= 0;
	where_in_block <= 0;
	
	data_in <= 8'd0;
	

end

always
begin
	#1 clk <= ~clk;
end

//inital reset and setup
always
begin
	//reset
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	//end reset and assert vld_crc
	@(posedge clk) begin
		reset <= 1'b0;
		vld_crc <= 1'b1;
	end
	//send code block size, start sending data
	@(posedge clk) begin
		vld_crc <= 1'b0;
		cbs <= 1'b0;
		start_rec <= 1'b1;
		counter <= 0;
		rdy_out <= 1'b1;
	end
	//wait until we get vld_out
	@(posedge vld_out) begin
		start_rec <= 1'b0;
	end
	@(posedge clk) begin
		rdy_out <= 1'b0;
		start_send <= 1'b1;
		counter <= 0;
	end
	#300
	$stop;
end

always @(posedge clk)
begin
	if(start_rec) begin
		$display("count: %0d | where: %0d | data_in: %b", counter, where_in_block, data_in);
		where_in_block = counter*8;	
		data_in = in[where_in_block +: 8];
		counter = counter+1;	
	end
	if(start_send) begin
		$display("count: %0d | where: %0d | data_out: %b | expected: %b | correct: %s", counter, where_in_block, data_out, expected_out[where_in_block +: 8], correct);
		where_in_block = counter*8;
		out[where_in_block +: 8] = data_out;
		if(out[where_in_block +: 8] == expected_out[where_in_block +: 8])
		begin
			correct = "TRUE";
		end
		else 
		begin
			correct = "FALSE";
		end
		counter = counter + 1;
	end
end

interleaver dut(clk, reset, vld_crc, rdy_out, cbs, data_in, rdy_crc, vld_out, data_out);


endmodule


